netcdf netcdf_simpleparticletest {
dimensions:
	time = UNLIMITED ;
	particleno = 3 ;
variables:
	float time(time);
	int particleno(time, particleno) ;
	float xpos(time, particleno) ;
	float ypos(time, particleno) ;
//	float xvel(time, particleno) ;
//	float yvel(time, particleno) ;
//	float pressure(time, particleno) ;
//	float density(time, particleno) ;
//	float depth(time, particleno) ;
data:

// data =
//  0, 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11,
//  12, 13, 14, 15, 16, 17, 18, 19, 20, 21, 22, 23,
//  24, 25, 26, 27, 28, 29, 30, 31, 32, 33, 34, 35,
//  36, 37, 38, 39, 40, 41, 42, 43, 44, 45, 46, 47,
//  48, 49, 50, 51, 52, 53, 54, 55, 56, 57, 58, 59,
//  60, 61, 62, 63, 64, 65, 66, 67, 68, 69, 70, 71 ;
	
	time = 1.01,2.01,3.01;
	particleno = 1,2,3,
	1,2,3,
	1,3,2;
	 xpos = 1,2,1.01,
	1,2,1.01,
	1,2,3.01;
	ypos = 0.0,0.0,0.01,
	0,0,0.02,
	0,0,0.03;
//	float xvel(particleno, time) ;
//	float yvel(particleno, time) ;
//	float pressure(particleno, time) ;
//	float density(particleno, time) ;
//	float depth(particleno, time) ;
}
